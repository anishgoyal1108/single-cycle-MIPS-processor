LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY PC IS
	PORT (
		clock : IN STD_LOGIC;
		PCin : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		PCout : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END PC;

ARCHITECTURE internal OF PC IS
	SIGNAL count : STD_LOGIC; 
BEGIN
	PROCESS (clock, PCin)
	BEGIN
		IF clock'EVENT AND clock = '1' THEN
			PCout <= PCin;
		END IF;
	END PROCESS;

END internal;