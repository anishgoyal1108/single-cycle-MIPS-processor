LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY Sign_Ext IS
	PORT (
		A : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		Y : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END Sign_Ext;

ARCHITECTURE internal OF Sign_Ext IS
BEGIN
	PROCESS (A)
	BEGIN
		IF a(15) = '0' THEN
			Y <= "0000000000000000" & A; 
		ELSIF a(15) = '1' THEN
			Y <= "1111111111111111" & A; 
		END IF; 
	END PROCESS;
END internal;