LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ShiftL2 IS
	PORT (
		A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Y : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END ShiftL2;

ARCHITECTURE internal OF ShiftL2 IS
BEGIN
	Y <= A(29 DOWNTO 0) & "00";
END internal;