LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY Adder IS
	PORT (
		x1, x2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Y : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END Adder;

ARCHITECTURE structure OF Adder IS
BEGIN
	Y <= x1 + x2;
END structure;